`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:36:39 11/06/2014 
// Design Name: 
// Module Name:    ROM_Seg 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ROM_Seg(
    input clk,
    input [3:0] dir,
    output reg[29:0] dato
	);

always@(posedge clk)
    case(dir)
   	 4'b0000: dato<= 30'b001011100010001011100010010001;
   	 4'b0001: dato<= 30'b010011100010011100010011100100;
   	 4'b0010: dato<= 30'b011001011011001011001011011001;
   	 4'b0011: dato<= 30'b011010010110001001010100011100;
   	 4'b0100: dato<= 30'b010100010010011100010001100011;
   	 4'b0101: dato<= 30'b001100001011010011001010001100;
   	 4'b0110: dato<= 30'b010011001010100001010001100010;
   	 4'b0111: dato<= 30'b100011010001010011010101100001;
   	 4'b1000: dato<= 30'b001010100001011010100011001100;
   	 4'b1001: dato<= 30'b100011010011010100001011001010;
   	 4'b1010: dato<= 30'b001100011010001010011100010100;
   	 4'b1011: dato<= 30'b100010001011100010001010100011;
   	 4'b1100: dato<= 30'b010100001010011100010011100001;
   	 4'b1101: dato<= 30'b001100011001010100011010001010;
   	 4'b1110: dato<= 30'b001001100011011010100001010011;
   	 4'b1111: dato<= 30'b001011001011001011001011001011;
    endcase

endmodule
